//-----------------------------------------------------------------
//                      Baseline JPEG Decoder
//                             V0.1
//                       Ultra-Embedded.com
//                        Copyright 2020
//
//                   admin@ultra-embedded.com
//-----------------------------------------------------------------
//                      License: Apache 2.0
// This IP can be freely used in commercial projects, however you may
// want access to unreleased materials such as verification environments,
// or test vectors, as well as changes to the IP for integration purposes.
// If this is the case, contact the above address.
// I am interested to hear how and where this IP is used, so please get
// in touch!
//-----------------------------------------------------------------
// Copyright 2020 Ultra-Embedded.com
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//-----------------------------------------------------------------


//Candidate for BSGMEM
module jpeg_idct_ram_dp
(
    // Inputs
     input           clk_i
    ,input           rst_i
    ,input  [  5:0]  addr0_i
    ,input  [ 15:0]  data0_i
    ,input           wr0_i
    // ,input           clk1_i
    // ,input           rst1_i
    ,input  [  5:0]  addr1_i
    ,input  [ 15:0]  data1_i
    ,input           wr1_i

    // Outputs
    ,output [ 15:0]  data0_o
    ,output [ 15:0]  data1_o
);



//-----------------------------------------------------------------
// Dual Port RAM
// Mode: Read First
//-----------------------------------------------------------------
/* verilator lint_off MULTIDRIVEN */
    //-----------------------------------------------------------------
    // LUT for decode values
    bsg_mem_1rw_sync #(.width_p(16)
                          , .els_p(64)
) jpeg_idct_ram_dp_mem1
   (.clk_i(clk_i)
    ,.reset_i(rst_i)
    ,.data_i(data0_i)
    ,.addr_i(addr0_i)
    , .v_i(1'b1)
    , .w_i(wr0_i)
    , .data_o(data0_o)
    );

        bsg_mem_1rw_sync #(.width_p(16)
                          , .els_p(64)
) jpeg_idct_ram_dp_mem2
   (.clk_i(clk_i)
    ,.reset_i(rst_i)
    ,.data_i(data1_i)
    ,.addr_i(addr1_i)
    , .v_i(1'b1)
    , .w_i(wr1_i)
    , .data_o(data1_o)
    );

// bsg_mem_2rw_sync #(.width_p(16)
//                            , .els_p(64)

// ) jpeg_idct_ram_dp_mem
//    (.clk_i(clk_i)
//     , .reset_i(rst_i)

//     , .a_v_i(1'b1)
//     , .a_addr_i(addr0_i)
//     , .a_data_i(data0_i)
//     ,.a_w_i(wr0_i)
//     , .b_v_i(1'b1)
//     , .b_addr_i(addr1_i)
//     , .b_data_i(data1_i)
//     ,.b_w_i(wr1_i)

//     // currently unused
//     , .a_data_o(data0_o)
//     , .b_data_o(data1_o)
//     );
// reg [15:0]   ram [63:0] /*verilator public*/;
// /* verilator lint_on MULTIDRIVEN */


// reg [15:0] ram_read0_q;
// reg [15:0] ram_read1_q;


// // Synchronous write
// always @ (posedge clk0_i)
// begin
//     if (wr0_i)
//         ram[addr0_i][15:0] <= data0_i[15:0];

//     ram_read0_q <= ram[addr0_i];
// end

// always @ (posedge clk1_i)
// begin
//     if (wr1_i)
//         ram[addr1_i][15:0] <= data1_i[15:0];

//     ram_read1_q <= ram[addr1_i];
// end


// assign data0_o = ram_read0_q;
// assign data1_o = ram_read1_q;

endmodule